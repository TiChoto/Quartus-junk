`timescale 1ns/1ps
module encoder_8to3_tb();
    reg [7:0] in;
    wire [2:0] out;
    
    encoder_8to3 inst (
	 .in(in), 
	 .out(out)
	 );
    
    initial begin
        $dumpfile("encoder_wave.vcd");
        $dumpvars(0, encoder_8to3_tb);
        
        #10 in = 8'b00000001; 
        #10 in = 8'b00000010; 
        #10 in = 8'b00000100; 
        #10 in = 8'b00001000; 
        #10 in = 8'b00010000; 
        #10 in = 8'b00100000;
        #10 in = 8'b01000000; 
        #10 in = 8'b10000000; 
        
    
        #10 in = 8'b00010010; 
        #10 in = 8'b00100100; 
        #10 in = 8'b11000000; 
        
        $finish;
    end
endmodule